11111            Waldo

11110000
11000011_11100011_00000001_11110000

11000011 11100011   
    1111 1


00111110       1
01111110       2	overlap question